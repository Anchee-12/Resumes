LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY REG IS
 PORT(GATE:IN STD_LOGIC;
      CLK:IN STD_LOGIC;
      DIN: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      DOUT:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END REG;
ARCHITECTURE BEHAV OF REG IS
BEGIN
 PROCESS(GATE,DIN)
 BEGIN
  IF CLK'EVENT AND CLK='1' THEN
   IF GATE='1' THEN DOUT<=DIN;
   END IF;
  END IF;
 END PROCESS;
END BEHAV;